test test test 
test test test
test test test 
